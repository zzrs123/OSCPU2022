module double_control(
    input a,
    input b,
    output f
);
  assign f = a ^ b;
endmodule
