// lab7的顶层模块 ps2_control
module ps2_control(

)